// Create a module that implements a NOT gate.

module top_module( inout in , output out);

  assign out = ~in;

endmodule